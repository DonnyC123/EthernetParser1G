package ddr_sdr_converter_pkg;

  typedef enum int {
    IDLE, 
    UPPER_HALF,
    LOWER_HALF
  } converter_state_t;

endpackage 