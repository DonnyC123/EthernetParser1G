package hash_table_pkg ();
  typedef enum logic {
    INSERT_QUERY  = 0,
    LOOK_UP_QUERY = 1
  } hash_query_t;

endpackage