package error_pulse_pkg;

  typedef enum logic {  
    NO_ERROR,
    ERROR
  } error_state_t;

endpackage